Since astronomers confirmed the presence of planets beyond our solar system, called exoplanets, humanity has wondered how many could harbor life. Now, we're one step closer to finding an answer. According to new research using data from NASA's retired planet-hunting mission, the Kepler space telescope, about half the stars similar in temperature to our Sun could have a rocky planet capable of supporting liquid water on its surface.

Our galaxy holds at least an estimated 300 million of these potentially habitable worlds, based on even the most conservative interpretation of the results in a new study to be published in The Astronomical Journal. Some of these exoplanets could even be our interstellar neighbors, with at least four potentially within 30 light-years of our Sun and the closest likely to be at most about 20 light-years from us. These are the minimum numbers of such planets based on the most conservative estimate that 7% of Sun-like stars host such worlds. However, at the average expected rate of 50%, there could be many more.

This research helps us understand the potential for these planets to have the elements to support life. This is an essential part of astrobiology, the study of life's origins and future in our universe.

The study is authored by NASA scientists who worked on the Kepler mission alongside collaborators from around the world. NASA retired the space telescope in 2018 after it ran out of fuel. Nine years of the telescope's observations revealed that there are billions of planets in our galaxy -- more planets than stars.

"Kepler already told us there were billions of planets, but now we know a good chunk of those planets might be rocky and habitable," said the lead author Steve Bryson, a researcher at NASA's Ames Research Center in California's Silicon Valley. "Though this result is far from a final value, and water on a planet's surface is only one of many factors to support life, it's extremely exciting that we calculated these worlds are this common with such high confidence and precision."

For the purposes of calculating this occurrence rate, the team looked at exoplanets between a radius of 0.5 and 1.5 times that of Earth's, narrowing in on planets that are most likely rocky. They also focused on stars similar to our Sun in age and temperature, plus or minus up to 1,500 degrees Fahrenheit.

That's a wide range of different stars, each with its own particular properties impacting whether the rocky planets in its orbit are capable of supporting liquid water. These complexities are partly why it is so difficult to calculate how many potentially habitable planets are out there, especially when even our most powerful telescopes can just barely detect these small planets. That's why the research team took a new approach.

Rethinking How to Identify Habitability

This new finding is a significant step forward in Kepler's original mission to understand how many potentially habitable worlds exist in our galaxy. Previous estimates of the frequency, also known as the occurrence rate, of such planets ignored the relationship between the star's temperature and the kinds of light given off by the star and absorbed by the planet.

The new analysis accounts for these relationships, and provides a more complete understanding of whether or not a given planet might be capable of supporting liquid water, and potentially life. That approach is made possible by combining Kepler's final dataset of planetary signals with data about each star's energy output from an extensive trove of data from the European Space Agency's Gaia mission.

"We always knew defining habitability simply in terms of a planet's physical distance from a star, so that it's not too hot or cold, left us making a lot of assumptions," said Ravi Kopparapu, an author on the paper and a scientist at NASA's Goddard Space Flight Center in Greenbelt, Maryland. "Gaia's data on stars allowed us to look at these planets and their stars in an entirely new way."

Gaia provided information about the amount of energy that falls on a planet from its host star based on a star's flux, or the total amount of energy that is emitted in a certain area over a certain time. This allowed the researchers to approach their analysis in a way that acknowledged the diversity of the stars and solar systems in our galaxy.

"Not every star is alike," said Kopparapu. "And neither is every planet."

Though the exact effect is still being researched, a planet's atmosphere figures into how much light is needed to allow liquid water on a planet's surface as well. Using a conservative estimate of the atmosphere's effect, the researchers estimated an occurrence rate of about 50% -- that is, about half of Sun-like stars have rocky planets capable of hosting liquid water on their surfaces. An alternative optimistic definition of the habitable zone estimates about 75%.

Kepler's Legacy Charts Future Research

This result builds upon a long legacy of work of analyzing Kepler data to obtain an occurrence rate and sets the stage for future exoplanet observations informed by how common we now expect these rocky, potentially habitable worlds to be. Future research will continue to refine the rate, informing the likelihood of finding these kinds of planets and feeding into plans for the next stages of exoplanet research, including future telescopes.

"Knowing how common different kinds of planets are is extremely valuable for the design of upcoming exoplanet-finding missions," said co-author Michelle Kunimoto, who worked on this paper after finishing her doctorate on exoplanet occurrence rates at the University of British Columbia, and recently joined the Transiting Exoplanet Survey Satellite, or TESS, team at the Massachusetts Institute of Technology in Cambridge, Massachusetts. "Surveys aimed at small, potentially habitable planets around Sun-like stars will depend on results like these to maximize their chance of success."

After revealing more than 2,800 confirmed planets outside our solar system, the data collected by the Kepler space telescope continues to yield important new discoveries about our place in the universe. Though Kepler's field of view covered only 0.25% of the sky, the area that would be covered by your hand if you held it up at arm's length towards the sky, its data has allowed scientists to extrapolate what the mission's data means for the rest of the galaxy. That work continues with TESS, NASA's current planet hunting telescope.

"To me, this result is an example of how much we've been able to discover just with that small glimpse beyond our solar system," said Bryson. "What we see is that our galaxy is a fascinating one, with fascinating worlds, and some that may not be too different from our own."